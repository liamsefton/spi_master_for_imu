module spi_master (
    input i_clk12,    //12 mhz system clk
    input i_rst,      //not really sure how to use resets yet

    input i_start_cmd,
    input i_rw_cmd,
    input [6:0] i_reg_addr,  //will be concatenated with i_rw_cmd to form the full address (with the rw bit being the most significant bit)
    input [7:0] i_wr_data,
    output reg [7:0] o_rd_data,
    output reg o_busy,

    output reg sclk,
    output reg mosi,
    output reg cs,     //active low (activate by setting low at start and deactivate at the end)
    input miso
);

localparam [1:0] IDLE = 2'b00;
localparam [1:0] SEND_ADDR = 2'b01;
localparam [1:0] DATA_HANDLER = 2'b10;
localparam [1:0] WAIT_CS = 2'b11;

localparam [4:0] CLK_DIV1 = 5'd12;  //rising edge amount for sclk
localparam [4:0] CLK_DIV2 = 5'd24;  //falling edge amount for sclk

reg sclk_rise, sclk_fall;    //generated by first state machine
reg [2:0] curr_state;

reg rw_cmd;  //0: write - 1: read

reg [6:0] reg_addr;
reg sclk_en;          //enables the slower clock for spi
reg [7:0] data_sreg;  //data_sreg no idea why this is needed

reg [4:0] clk_cnt = 5'b00000;     //this is the system clock counter that generates the rising and falling edges of sclk

always @(posedge i_clk12 or posedge i_rst)
begin
    if(i_rst)
    begin
        clk_cnt <= 5'b00000;
        sclk_rise <= 1'b0;
        sclk_fall <= 1'b0;
        sclk <= 1'b1;  //changed to reflect imu datasheet
    end
    else
    begin
        sclk_rise <= 1'b0;
        sclk_fall <= 1'b0;

        if(sclk_en)
        begin
            clk_cnt <= clk_cnt + 1;
            if(clk_cnt == CLK_DIV1)
            begin
                sclk_rise <= 1'b1;
                sclk <= 1'b1;
            end
            if(clk_cnt == CLK_DIV2)
            begin
                sclk_fall <= 1'b1;
                sclk <= 1'b0;
                clk_cnt = 5'b00000;
            end
        end
        else
        begin
            clk_cnt <= 5'b00000;
            sclk <= 1'b1;  //changed to reflect imu datasheet
        end
    end
end

reg [1:0] bit_cnt;

always @(posedge i_clk12 or posedge i_rst)
begin
    if(i_rst)
    begin
        o_busy <= 1'b0;
        o_rd_data <= 8'h00;
        sclk_en <= 1'b0;
        mosi <= 1'b0;
        bit_cnt <= 3'b000;
        rw_cmd <= 1'b0;
        reg_addr <= 7'h0;
        data_sreg <= 8'h00;
        curr_state <= IDLE;
        cs <= 1'b1;
    end
    else
    begin
        case(curr_state)
            IDLE:
            begin
                o_busy <= 1'b0;
                cs <= 1'b1;
                mosi <= 1'b0;
                sclk_en <= 1'b0;
                bit_cnt <= 4'h0;
                rw_cmd <= 1'b0;
                reg_addr <= 7'h0;
                data_sreg <= 8'h00;

                if(i_start_cmd)
                begin
                    if(!i_rw_cmd)
                    begin
                        rw_cmd <= 1'b0;
                        data_sreg <= i_wr_data;
                    end
                    else //read
                    begin
                        rw_cmd <= 1'b1;
                        data_sreg <= 8'h00;
                    end

                    o_busy <= 1'b1;
                    cs <= 1'b0;
                    sclk_en <= 1'b1;
                    reg_addr <= i_reg_addr;
                    curr_state <= SEND_ADDR;
                end
            end
            SEND_ADDR:
            begin
                if(sclk_fall)
                begin
                    if(bit_cnt == 3'b000)
                    begin
                        mosi <= rw_cmd;
                    end
                    else
                    begin
                        mosi <= reg_addr[7-bit_cnt];
                    end
                    if(bit_cnt == 3'd7)
                    begin
                        bit_cnt <= 3'h0;
                        curr_state <= DATA_HANDLER;
                    end
                    else
                    begin
                        bit_cnt <= bit_cnt + 1;
                    end
                end
            end
            DATA_HANDLER:
            begin
                if(sclk_rise)
                begin
                    if(rw_cmd)
                    begin
                        data_sreg[0] <= miso;
                        data_sreg[7:1] <= data_sreg[6:0];
                    end
                end
                if(sclk_fall)
                begin
                    if(!rw_cmd)
                    begin
                        mosi <= data_sreg[7-bit_cnt];
                    end
                    if(bit_cnt == 3'd7)
                    begin
                        bit_cnt <= 3'd0;
                        if(rw_cmd)
                        begin
                            o_rd_data <= data_sreg;
                        end
                        curr_state <= WAIT_CS;
                    end
                    else
                    begin
                        bit_cnt <= bit_cnt + 1;
                    end
                end
            end
            WAIT_CS:
            begin
                if(bit_cnt == 3'd7)
                begin
                    cs <= 1'b1;
                    sclk_en <= 1'b0;
                    o_busy <= 1'b0;
                    mosi <= 1'b0;
                    curr_state <= IDLE;
                    bit_cnt <= 0;
                end
                else
                begin
                    bit_cnt <= bit_cnt + 1;
                end
            end
        endcase
    end
end

endmodule



